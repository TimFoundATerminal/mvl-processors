module control(clock, 
    opcode, is_alu_operation,
    do_fetch, do_load, do_alu, do_mem_load, do_mem_store, do_reg_store, do_next, do_reset, do_halt,
    state);

    /* 
    Control Module for the CPU

    Does not need to take any signals from a Bus as this system does not have any I/O devices
    */

    `include "parameters.vh"

    input wire clock;

    input wire [OPCODE_SIZE-1:0] opcode;
    input wire is_alu_operation;

    output wire do_fetch, do_load, do_alu, do_mem_load, do_mem_store, do_reg_store, do_next, do_reset, do_halt;

    output reg [3:0] state = `STATE_INSMEM_LOAD;

    always @(posedge clock) begin
        $display("State: %d, Opcode: %d", state, opcode);

        case (state)
            `STATE_RESET: begin
                state <= `STATE_FETCH;
            end

            `STATE_FETCH: begin
                state <= `STATE_REGLOAD;
            end

            `STATE_REGLOAD: begin
                if (is_alu_operation) 
                    state <= `STATE_ALU;
                else case (opcode)
                    // TODO MV operation
                    `LOAD:
                        state <= `STATE_LOAD;
                    `STORE:
                        state <= `STATE_STORE;
                    `LUI:
                        state <= `STATE_REGSTORE;
                    `LI:
                        state <= `STATE_REGSTORE;
                    `BEQ:
                        state <= `STATE_NEXT;
                    `BNE:
                        state <= `STATE_NEXT;
                    `HALT:
                        state <= `STATE_HALT;
                endcase
            end

            `STATE_ALU: begin
                state <= `STATE_REGSTORE;
            end

            `STATE_REGSTORE: begin
                state <= `STATE_NEXT;
            end

            `STATE_LOAD: begin
                state <= `STATE_REGSTORE;
            end

            `STATE_STORE: begin
                state <= `STATE_NEXT;
            end

            `STATE_NEXT: begin
                state <= `STATE_FETCH;
            end

            // explicit declaration of halt state
            `STATE_HALT: begin
                state <= `STATE_HALT;
            end

        endcase
    end

    // Control the CPU with the following signals
    assign do_fetch = (state == `STATE_FETCH);
    assign do_load = (state == `STATE_REGLOAD);
    assign do_alu = (state == `STATE_ALU);
    assign do_mem_load = (state == `STATE_LOAD);
    assign do_mem_store = (state == `STATE_STORE);
    assign do_reg_store = (state == `STATE_REGSTORE);
    assign do_next = (state == `STATE_NEXT);
    assign do_reset = (state == `STATE_RESET);
    assign do_halt = (state == `STATE_HALT);

endmodule