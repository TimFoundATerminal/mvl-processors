package ternary_package;
    parameter VPOS = 5.0;
    parameter VZERO = 0.0;
    parameter VNEG = -5.0;
    parameter VTHRESH_POS = 2.5;
    parameter VTHRESH_NEG = -2.5;
    parameter VDD = 5.0;
    parameter VSS = -5.0;
endpackage